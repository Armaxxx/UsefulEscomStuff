library ieee;
use ieee.std_logic_1164.all;
library lattice;
use lattice.all;
use packagemult4bit00.all;

entity topmult4bit00 is
  port(
       Am: in std_logic_vector(3 downto 0);
	   Bm: in std_logic_vector(3 downto 0);
       Rm: out std_logic_vector(7 downto 0));
end topmult4bit00;

architecture topmult4bit0 of topmult4bit00 is
signal S1, S2, S4: std_logic_vector(3 downto 0);
signal S5, S7, S8: std_logic_vector(3 downto 0);
signal S0, S3, S6: std_logic_vector(2 downto 0);
begin

  M00: and00 port map(Aa => Am(0),
                      Ba => Bm(0),
                      Ya => Rm(0));
  
  M01: and00 port map(Aa => Am(1),
                      Ba => Bm(0),
                      Ya => S0(0));
  
  M02: and00 port map(Aa => Am(2),
                      Ba => Bm(0),
                      Ya => S0(1));
  
  M03: and00 port map(Aa => Am(3),
                      Ba => Bm(0),
                      Ya => S0(2));

  M04: and00 port map(Aa => Am(0),
                      Ba => Bm(1),
                      Ya => S1(0));

  M05: and00 port map(Aa => Am(1),
                      Ba => Bm(1),
                      Ya => S1(1));

  M06: and00 port map(Aa => Am(2),
                      Ba => Bm(1),
                      Ya => S1(2));

  M07: and00 port map(Aa => Am(3),
                      Ba => Bm(1),
                      Ya => S1(3));

  M08: fa00 port map(C00 => '0',
                     A00 => S0(0),
					 B00 => S1(0),
					 C01 => S2(0),
                     S00 => Rm(1));
  
  M09: fa00 port map(C00 => S2(0),
                     A00 => S0(1),
					 B00 => S1(1),
					 C01 => S2(1),
                     S00 => S3(0));

  
  M10: fa00 port map(C00 => S2(1),
                     A00 => S0(2),
					 B00 => S1(2),
					 C01 => S2(2),
                     S00 => S3(1));
  
  M11: fa00 port map(C00 => S2(2),
                     A00 => '0',
					 B00 => S1(3),
					 C01 => S2(3),
                     S00 => S3(2));
					 
  M12: and00 port map(Aa => Am(0),
                      Ba => Bm(2),
                      Ya => S4(0));

  M13: and00 port map(Aa => Am(1),
                      Ba => Bm(2),
                      Ya => S4(1));

  M14: and00 port map(Aa => Am(2),
                      Ba => Bm(2),
                      Ya => S4(2));

  M15: and00 port map(Aa => Am(3),
                      Ba => Bm(2),
                      Ya => S4(3));

  M16: fa00 port map(C00 => '0',
                     A00 => S3(0),
                     B00 => S4(0),
					 C01 => S5(0),
                     S00 => Rm(2));

  M17: fa00 port map(C00 => S5(0),
                     A00 => S3(1),
                     B00 => S4(1),
					 C01 => S5(1),
                     S00 => S6(0));

  M18: fa00 port map(C00 => S5(1),
                     A00 => S3(2),
                     B00 => S4(2),
					 C01 => S5(2),
                     S00 => S6(1));


  M19: fa00 port map(C00 => S5(2),
                     A00 => S2(3),
                     B00 => S4(3),
					 C01 => S5(3),
                     S00 => S6(2));

  M20: and00 port map(Aa => Am(0),
                      Ba => Bm(3),
                      Ya => S7(0));

  M21: and00 port map(Aa => Am(1),
                      Ba => Bm(3),
                      Ya => S7(1));

  M22: and00 port map(Aa => Am(2),
                      Ba => Bm(3),
                      Ya => S7(2));

  M23: and00 port map(Aa => Am(3),
                      Ba => Bm(3),
                      Ya => S7(3));

  M24: fa00 port map(C00 => '0',
                     A00 => S6(0),
					 B00 => S7(0),
					 C01 => S8(0),
                     S00 => Rm(3));

  M25: fa00 port map(C00 => S8(0),
                     A00 => S6(1),
					 B00 => S7(1),
					 C01 => S8(1),
                     S00 => Rm(4));

  M26: fa00 port map(C00 => S8(1),
                     A00 => S6(2),
					 B00 => S7(2),
					 C01 => S8(2),
                     S00 => Rm(5));
					 
  M27: fa00 port map(C00 => S8(2),
                     A00 => S5(3),
					 B00 => S7(3),
					 C01 => Rm(7),
                     S00 => Rm(6));

end topmult4bit0;